package BlueXLNX;

import BSCANE2 :: *;
import BUFG :: *;
import BUFGCE :: *;
import GLBL :: *;
import IBUFDS :: *;
import JTAG_SIME2 :: *;
import MMCME4_ADV :: *;
import DiffClockAdapter :: *;

export BSCANE2 :: *;
export BUFG :: *;
export BUFGCE :: *;
export GLBL :: *;
export IBUFDS :: *;
export JTAG_SIME2 :: *;
export MMCME4_ADV :: *;
export DiffClockAdapter :: *;

endpackage